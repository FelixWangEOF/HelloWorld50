module hello;
    initial begin
        $display("hello world");
    end
endmodule 